`timescale 1ns/1ns

module caf_fpga(input sysclk);
endmodule // caf_fpga
